-------------------------------------------------------------------------------
-- Title      : Xilinx 7-series GTP Transceiver Tile
-- Project    : Open Communication Controller
-------------------------------------------------------------------------------
-- Author     : Daniel Tavares
-- Company    : CNPEM LNLS-DIG
-- Created    : 2020-04-30
-- Platform   : Xilinx
-------------------------------------------------------------------------------
-- Description: Encapsulates Xilinx 7-series GTP transceiver and corresponding
-- PLL and clock buffers with the settings required by the Open Communication
-- Controller protocol. One tile instance comprehends 1 to 4 transceivers.
--
-- Based on code generated by Vivado GT wizard (gtrxreset_seq.vhd) for the
-- receiver reset sequence (AR# 53561).
-------------------------------------------------------------------------------
--
-- Copyright (c) 2020 CNPEM
--
-- This source describes open hardware and is licensed under the CERN-OHL-W v2.
--
-- You may redistribute and modify this documentation and make products using
-- it under the terms of the CERN-OHL-W v2 (https:/cern.ch/cern-ohl, or (at
-- your option) any later version. This documentation is distributed WITHOUT
-- ANY EXPRESS OR IMPLIED WARRANTY, INCLUDING OF MERCHANTABILITY, SATISFACTORY
-- QUALITY AND FITNESS FOR A PARTICULAR PURPOSE. Please see the CERN-OHL-W v2
-- for applicable conditions.
--
-------------------------------------------------------------------------------

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

library unisim;
use unisim.vcomponents.all;

entity occ_gtpe2_tile is
generic
(
  g_SIMULATION            : string  := "FALSE";
  g_SIMULATION_SPEEDUP    : string  := "FALSE";
  g_NUM_CHANNELS          : integer range 1 to 4 := 1;  -- TODO: g_NUM_CHANNELS should range from 1 to 4
  g_REFCLK                : string  := "REFCLK0";       -- TODO: select among "REFCLK0", "REFCLK1", "EASTREFCLK0", "EASTREFCLK1", "WESTREFCLK0", "WESTREFCLK1"
  g_PHYSICAL_LAYER        : string  := "SFP"
);
port
(
  -----------------
  -- EXTERNAL PADS
  -----------------
  rxn_i                   : in  std_logic;
  rxp_i                   : in  std_logic;
  txn_o                   : out std_logic;
  txp_o                   : out std_logic;

  -----------------
  -- RECEIVER (RX)
  -----------------
  -- Reset
  rxreset_i               : in  std_logic;
  rxresetdone_o           : out std_logic;
  -- 8b10b Decoder
  rxcharisk_o             : out std_logic_vector(1 downto 0);
  rxdisperr_o             : out std_logic_vector(1 downto 0);
  rxnotintable_o          : out std_logic_vector(1 downto 0);
  -- Comma Detection and Alignment
  rxbyteisaligned_o       : out std_logic;
  rxbyterealign_o         : out std_logic;
  rxencommaalign_i        : in  std_logic;
  -- Elastic Buffer
  rxbufstatus_o           : out std_logic_vector(2 downto 0);
  -- Data Path Interface
  rxdata_o                : out std_logic_vector(15 downto 0);
  rxuserrdy_i             : in  std_logic;

  --------------------
  -- TRANSMITTER (TX)
  --------------------
  -- Reset
  txreset_i               : in  std_logic;
  txresetdone_o           : out std_logic;
  -- 8b10b Encoder
  txcharisk_i             : in  std_logic_vector(1 downto 0);
  -- Data Path Interface
  txdata_i                : in  std_logic_vector(15 downto 0);
  txuserrdy_i             : in  std_logic;

  -------------
  -- GT CLOCKS
  -------------
  -- Input clocks
  refclk0_i               : in std_logic;
  refclk1_i               : in std_logic;

  -- Output clocks to be used by user logic
  usrclk_o                : out std_logic;

  -----------------------
  -- RX/TX CONFIGURATION
  -----------------------
  loopback_i              : in  std_logic_vector(2 downto 0);
  powerdown_i             : in  std_logic_vector(1 downto 0);

  -------
  -- PLL
  -------
  -- Clock for PLL lock detection circuit
  pll_lockdetclk_i        : in  std_logic;
  pll_lock_o              : out std_logic;
  pll_refclklost_o        : out std_logic;
  pll_refclksel_i         : in  std_logic_vector(2 downto 0);
  pll_rst_i               : in  std_logic;
  
  ------------------
  -- INITIALIZATION
  ------------------
  -- Used on reset sequence workaround (AR# 53561)
  init_rst_i              : in  std_logic;
  init_clk_i              : in  std_logic
);
end occ_gtpe2_tile;

architecture rtl of occ_gtpe2_tile is

  -- PLL dividers configuration
  constant c_PLLFBDIV       : integer := 5;
  constant c_PLLFBDIV45     : integer := 5;
  constant c_PLLREFDIV      : integer := 1;

  -- Clock signals
  signal usrclk             : std_logic;
  signal txoutclk           : std_logic;
  signal pll0clk            : std_logic;
  signal pll0refclk         : std_logic;
  signal pll1clk            : std_logic;
  signal pll1refclk         : std_logic;

  -- Datapath signals
  signal rxdata             : std_logic_vector(31 downto 0);
  signal txdata             : std_logic_vector(31 downto 0);
  signal rxcharisk          : std_logic_vector(3 downto 0);
  signal rxdisperr          : std_logic_vector(3 downto 0);
  signal rxnotintable       : std_logic_vector(3 downto 0);

  -- RX reset sequence signals (AR# 53561)
  signal rxpmaresetdone     : std_logic;
  signal txpmaresetdone     : std_logic;
  signal rxreset            : std_logic;
  signal drp_op_done        : std_logic;
  signal drpaddr            : std_logic_vector(8 downto 0);
  signal drpen              : std_logic;
  signal drpwe              : std_logic;
  signal drpdo              : std_logic_vector(15 downto 0);
  signal drpdi              : std_logic_vector(15 downto 0);
  signal drprdy             : std_logic;

  -- RX reset sequence component (AR# 53561)
  component gtrxreset_seq_sim
  port ( 
    RST             : in  std_logic;
    GTRXRESET_IN    : in  std_logic;
    RXPMARESETDONE  : in  std_logic;
    GTRXRESET_OUT   : out std_logic;  
    DRPCLK          : in  std_logic;
    DRPADDR         : out std_logic_vector(8 downto 0);
    DRPDO           : in  std_logic_vector(15 downto 0);
    DRPDI           : out std_logic_vector(15 downto 0);
    DRPRDY          : in  std_logic;
    DRPEN           : out std_logic;
    DRPWE           : out std_logic;
    DRP_OP_DONE     : out std_logic
  );
  end component;

  component gtrxreset_seq
  port ( 
    RST             : in  std_logic;
    GTRXRESET_IN    : in  std_logic;
    RXPMARESETDONE  : in  std_logic;
    GTRXRESET_OUT   : out std_logic;  
    DRPCLK          : in  std_logic;
    DRPADDR         : out std_logic_vector(8 downto 0);
    DRPDO           : in  std_logic_vector(15 downto 0);
    DRPDI           : out std_logic_vector(15 downto 0);
    DRPRDY          : in  std_logic;
    DRPEN           : out std_logic;
    DRPWE           : out std_logic;
    DRP_OP_DONE     : out std_logic
  );
  end component;

begin

  -- Trim/pad data
  rxdata_o        <= rxdata(15 downto 0);
  txdata          <= "0000000000000000" & txdata_i;
  rxcharisk_o     <= rxcharisk(1 downto 0);
  rxdisperr_o     <= rxdisperr(1 downto 0);
  rxnotintable_o  <= rxnotintable(1 downto 0);

  -- GTPE2_CHANNEL instances
  cmp_gtpe2_0 : GTPE2_CHANNEL
  generic map
  (
    -- Simulation
    SIM_RECEIVER_DETECT_PASS        => "TRUE",
    SIM_RESET_SPEEDUP               => g_SIMULATION_SPEEDUP,
    SIM_TX_EIDLE_DRIVE_LEVEL        => "X",
    SIM_VERSION                     => "2.0",
    -- RX Byte and Word Alignment   
    ALIGN_COMMA_DOUBLE              => "FALSE",
    ALIGN_COMMA_ENABLE              => "1111111111",
    ALIGN_COMMA_WORD                => 1,
    ALIGN_MCOMMA_DET                => "TRUE",
    ALIGN_MCOMMA_VALUE              => "1010000011", -- -K28.5+ (10-bit symbol)
    ALIGN_PCOMMA_DET                => "TRUE",
    ALIGN_PCOMMA_VALUE              => "0101111100", -- +K28.5- (10-bit symbol)
    SHOW_REALIGN_COMMA              => "FALSE",
    RXSLIDE_AUTO_WAIT               => 7,
    RXSLIDE_MODE                    => "OFF", -- INFO: "PCS" for manual alignment
    RX_SIG_VALID_DLY                => 10,
    -- RX 8B/10B Decoder            
    RX_DISPERR_SEQ_MATCH            => "TRUE",
    DEC_MCOMMA_DETECT               => "TRUE",
    DEC_PCOMMA_DETECT               => "TRUE",
    DEC_VALID_COMMA_ONLY            => "FALSE",
    -- RX Clock Correction          
    CBCC_DATA_SOURCE_SEL            => "DECODED",
    CLK_COR_SEQ_2_USE               => "FALSE",
    CLK_COR_KEEP_IDLE               => "FALSE",
    CLK_COR_MAX_LAT                 => 15,    -- TODO: check if it can be improved (i.e. reduced)
    CLK_COR_MIN_LAT                 => 12,    -- TODO: check if it can be improved (i.e. reduced)
    CLK_COR_PRECEDENCE              => "TRUE",
    CLK_COR_REPEAT_WAIT             => 0,
    CLK_COR_SEQ_LEN                 => 2,
    CLK_COR_SEQ_1_ENABLE            => "1111",
    CLK_COR_SEQ_1_1                 => "0110111100", -- K28.5 (8-bit symbol)
    CLK_COR_SEQ_1_2                 => "0010010101", -- D21.4 (8-bit symbol)
    CLK_COR_SEQ_1_3                 => "0000000000",
    CLK_COR_SEQ_1_4                 => "0000000000",
    CLK_CORRECT_USE                 => "TRUE",
    CLK_COR_SEQ_2_ENABLE            => "1111",
    CLK_COR_SEQ_2_1                 => "0000000000",
    CLK_COR_SEQ_2_2                 => "0000000000",
    CLK_COR_SEQ_2_3                 => "0000000000",
    CLK_COR_SEQ_2_4                 => "0000000000",
    -- RX Channel Bonding           
    CHAN_BOND_KEEP_ALIGN            => "FALSE",
    CHAN_BOND_MAX_SKEW              => 1,
    CHAN_BOND_SEQ_LEN               => 1,
    CHAN_BOND_SEQ_1_1               => "0000000000",
    CHAN_BOND_SEQ_1_2               => "0000000000",
    CHAN_BOND_SEQ_1_3               => "0000000000",
    CHAN_BOND_SEQ_1_4               => "0000000000",
    CHAN_BOND_SEQ_1_ENABLE          => "1111",
    CHAN_BOND_SEQ_2_1               => "0000000000",
    CHAN_BOND_SEQ_2_2               => "0000000000",
    CHAN_BOND_SEQ_2_3               => "0000000000",
    CHAN_BOND_SEQ_2_4               => "0000000000",
    CHAN_BOND_SEQ_2_ENABLE          => "1111",
    CHAN_BOND_SEQ_2_USE             => "FALSE",
    FTS_DESKEW_SEQ_ENABLE           => "1111",
    FTS_LANE_DESKEW_CFG             => "1111",
    FTS_LANE_DESKEW_EN              => "FALSE",
    -- RX Margin Analysis           
    ES_CONTROL                      => "000000",
    ES_ERRDET_EN                    => "FALSE",
    ES_EYE_SCAN_EN                  => "FALSE",
    ES_HORZ_OFFSET                  => x"010",
    ES_PMA_CFG                      => "0000000000",
    ES_PRESCALE                     => "00000",
    ES_QUALIFIER                    => x"00000000000000000000",
    ES_QUAL_MASK                    => x"00000000000000000000",
    ES_SDATA_MASK                   => x"00000000000000000000",
    ES_VERT_OFFSET                  => "000000000",
    -- RX FPGA Interface            
    RX_DATA_WIDTH                   => 20,
    -- PMA                          
    OUTREFCLK_SEL_INV               => "11",
    PMA_RSV                         => x"00000333",
    PMA_RSV2                        => x"00002040",
    PMA_RSV3                        => "00",
    PMA_RSV4                        => "0000",
    RX_BIAS_CFG                     => "0000111100110011",
    DMONITOR_CFG                    => x"000A00",
    RX_CM_SEL                       => "01",   -- TODO: check physical interface
    RX_CM_TRIM                      => "0000", -- TODO: check physical interface / AFC-timing uses 1010
    RX_DEBUG_CFG                    => "00000000000000",
    RX_OS_CFG                       => "0000010000000",
    TERM_RCAL_CFG                   => "100001000010000",
    TERM_RCAL_OVRD                  => "000",
    TST_RSV                         => x"00000000",
    RX_CLK25_DIV                    => 5, -- TODO: operates for refclk up to 125 MHz only? Look at UG196
    TX_CLK25_DIV                    => 5, -- TODO: operates for refclk up to 125 MHz only? Look at UG196
    UCODEER_CLR                     => '0',
    -- PCI Express                  
    PCS_PCIE_EN                     => "FALSE",
    -- PCS                          
    PCS_RSVD_ATTR                   => x"000000000000",
    -- RX Buffer                    
    RXBUF_ADDR_MODE                 => "FULL",
    RXBUF_EIDLE_HI_CNT              => "1000",
    RXBUF_EIDLE_LO_CNT              => "0000",
    RXBUF_EN                        => "TRUE",
    RX_BUFFER_CFG                   => "000000",
    RXBUF_RESET_ON_CB_CHANGE        => "TRUE",
    RXBUF_RESET_ON_COMMAALIGN       => "FALSE",
    RXBUF_RESET_ON_EIDLE            => "FALSE",
    RXBUF_RESET_ON_RATE_CHANGE      => "TRUE",
    RXBUFRESET_TIME                 => "00001",
    RXBUF_THRESH_OVFLW              => 61,
    RXBUF_THRESH_OVRD               => "FALSE",
    RXBUF_THRESH_UNDFLW             => 4,
    RXDLY_CFG                       => x"001F",
    RXDLY_LCFG                      => x"030",
    RXDLY_TAP_CFG                   => x"0000",
    RXPH_CFG                        => x"C00002",
    RXPHDLY_CFG                     => x"084020",
    RXPH_MONITOR_SEL                => "00000",
    RX_XCLK_SEL                     => "RXREC",
    RX_DDI_SEL                      => "000000",
    RX_DEFER_RESET_BUF_EN           => "TRUE",
    -- CDR                          
    RXCDR_CFG                       => x"0000107FE406001041010",  -- INFO: depends on RXOUT_DIV attribute
    RXCDR_FR_RESET_ON_EIDLE         => '0',
    RXCDR_HOLD_DURING_EIDLE         => '0',
    RXCDR_PH_RESET_ON_EIDLE         => '0',
    RXCDR_LOCK_CFG                  => "001001",
    -- RX Initialization and Reset  
    RXCDRFREQRESET_TIME             => "00001",
    RXCDRPHRESET_TIME               => "00001",
    RXISCANRESET_TIME               => "00001",
    RXPCSRESET_TIME                 => "00001",
    RXPMARESET_TIME                 => "00011",
    -- RX OOB Signalling            
    RXOOB_CFG                       => "0000110",
    -- RX Gearbox                   
    RXGEARBOX_EN                    => "FALSE",
    GEARBOX_MODE                    => "000",
    -- PRBS Detection               
    RXPRBS_ERR_LOOPBACK             => '0',
    -- Power-Down                   
    PD_TRANS_TIME_FROM_P2           => x"03c",
    PD_TRANS_TIME_NONE_P2           => x"3c",
    PD_TRANS_TIME_TO_P2             => x"64",
    -- RX OOB Signalling            
    SAS_MAX_COM                     => 64,
    SAS_MIN_COM                     => 36,
    SATA_BURST_SEQ_LEN              => "0101",
    SATA_BURST_VAL                  => "100",
    SATA_EIDLE_VAL                  => "100",
    SATA_MAX_BURST                  => 8,
    SATA_MAX_INIT                   => 21,
    SATA_MAX_WAKE                   => 7,
    SATA_MIN_BURST                  => 4,
    SATA_MIN_INIT                   => 12,
    SATA_MIN_WAKE                   => 4,
    -- RX Fabric Clock Output Control
    TRANS_TIME_RATE                 => x"0E",
    -- TX Buffer                    
    TXBUF_EN                        => "TRUE",
    TXBUF_RESET_ON_RATE_CHANGE      => "TRUE",
    TXDLY_CFG                       => x"001F",
    TXDLY_LCFG                      => x"030",
    TXDLY_TAP_CFG                   => x"0000",
    TXPH_CFG                        => x"0780",
    TXPHDLY_CFG                     => x"084020",
    TXPH_MONITOR_SEL                => "00000",
    TX_XCLK_SEL                     => "TXOUT",
    -- TX FPGA Interface            
    TX_DATA_WIDTH                   => 20,
    -- TX Configurable Driver       
    TX_DEEMPH0                      => "000000",
    TX_DEEMPH1                      => "000000",
    TX_EIDLE_ASSERT_DELAY           => "110",
    TX_EIDLE_DEASSERT_DELAY         => "100",
    TX_LOOPBACK_DRIVE_HIZ           => "FALSE",
    TX_MAINCURSOR_SEL               => '0',
    TX_DRIVE_MODE                   => "DIRECT",
    TX_MARGIN_FULL_0                => "1001110",
    TX_MARGIN_FULL_1                => "1001001",
    TX_MARGIN_FULL_2                => "1000101",
    TX_MARGIN_FULL_3                => "1000010",
    TX_MARGIN_FULL_4                => "1000000",
    TX_MARGIN_LOW_0                 => "1000110",
    TX_MARGIN_LOW_1                 => "1000100",
    TX_MARGIN_LOW_2                 => "1000010",
    TX_MARGIN_LOW_3                 => "1000000",
    TX_MARGIN_LOW_4                 => "1000000",
    -- TX Gearbox                   
    TXGEARBOX_EN                    => "FALSE",
    -- TX Initialization and Reset  
    TXPCSRESET_TIME                 => "00001",
    TXPMARESET_TIME                 => "00001",
    -- TX Receiver Detection        
    TX_RXDETECT_CFG                 => x"1832",
    TX_RXDETECT_REF                 => "100",
    -- JTAG                         
    ACJTAG_DEBUG_MODE               => '0',
    ACJTAG_MODE                     => '0',
    ACJTAG_RESET                    => '0',
    -- CDR                          
    CFOK_CFG                        => x"49000040E80",
    CFOK_CFG2                       => "0100000",
    CFOK_CFG3                       => "0100000",
    CFOK_CFG4                       => '0',
    CFOK_CFG5                       => x"0",
    CFOK_CFG6                       => "0000",
    RXOSCALRESET_TIME               => "00011",
    RXOSCALRESET_TIMEOUT            => "00000",
    -- PMA                          
    CLK_COMMON_SWING                => '0',
    RX_CLKMUX_EN                    => '1',
    TX_CLKMUX_EN                    => '1',
    ES_CLK_PHASE_SEL                => '0',
    USE_PCS_CLK_PHASE_SEL           => '0',
    PMA_RSV6                        => '0',
    PMA_RSV7                        => '0',
    -- TX Configuration Driver      
    TX_PREDRIVER_MODE               => '0',
    PMA_RSV5                        => '0',
    SATA_PLL_CFG                    => "VCO_3000MHZ",
    -- RX Fabric Clock Output Control
    RXOUT_DIV                       => 1,   -- INFO: affects RXCDR_CFG attribute
    -- TX Fabric Clock Output Control
    TXOUT_DIV                       => 1,   -- INFO: affects RXCDR_CFG attribute
    -- RX Phase Interpolator
    RXPI_CFG0                       => "000",
    RXPI_CFG1                       => '1',
    RXPI_CFG2                       => '1',
    -- RX Equalizer
    ADAPT_CFG0                      => x"00000",
    RXLPMRESET_TIME                 => "0001111",
    RXLPM_BIAS_STARTUP_DISABLE      => '0',
    RXLPM_CFG                       => "0110",
    RXLPM_CFG1                      => '0',
    RXLPM_CM_CFG                    => '0',
    RXLPM_GC_CFG                    => "111100010",
    RXLPM_GC_CFG2                   => "001",
    RXLPM_HF_CFG                    => "00001111110000",
    RXLPM_HF_CFG2                   => "01010",
    RXLPM_HF_CFG3                   => "0000",
    RXLPM_HOLD_DURING_EIDLE         => '0',
    RXLPM_INCM_CFG                  => '0', -- TODO: check physical interface
    RXLPM_IPCM_CFG                  => '1', -- TODO: check physical interface
    RXLPM_LF_CFG                    => "000000001111110000",
    RXLPM_LF_CFG2                   => "01010",
    RXLPM_OSINT_CFG                 => "100",
    -- TX Phase Interpolator PPM Controller
    TXPI_CFG0                       => "00",
    TXPI_CFG1                       => "00",
    TXPI_CFG2                       => "00",
    TXPI_CFG3                       => '0',
    TXPI_CFG4                       => '0',
    TXPI_CFG5                       => "000",
    TXPI_GREY_SEL                   => '0',
    TXPI_INVSTROBE_SEL              => '0',
    TXPI_PPMCLK_SEL                 => "TXUSRCLK2",
    TXPI_PPM_CFG                    => x"00",
    TXPI_SYNFREQ_PPM                => "001", -- TODO: check this. Aurora and many other projects use 000, but gt wizard generated 001
    -- Loopback
    LOOPBACK_CFG                    => '0',
    PMA_LOOPBACK_CFG                => '0',
    -- RX OOB Signalling
    RXOOB_CLK_CFG                   => "PMA",
    -- TX OOB Signalling
    TXOOB_CFG                       => '0',
    -- RX Buffer
    RXSYNC_MULTILANE                => '0',
    RXSYNC_OVRD                     => '0',
    RXSYNC_SKIP_DA                  => '0',
    -- TX Buffer
    TXSYNC_MULTILANE                => '0',
    TXSYNC_OVRD                     => '0',
    TXSYNC_SKIP_DA                  => '0'
  )
  port map
  (
    -- CPLL
    GTRSVD                          => "0000000000000000",
    PCSRSVDIN                       => "0000000000000000",
    TSTIN                           => "11111111111111111111",
    -- Dynamic Reconfiguration Port (DRP)
    DRPADDR                         => drpaddr,
    DRPCLK                          => init_clk_i,
    DRPDI                           => drpdi,
    DRPDO                           => drpdo,
    DRPEN                           => drpen,
    DRPRDY                          => drprdy,
    DRPWE                           => drpwe,
    -- Clocking
    RXSYSCLKSEL                     => "00",   -- use PLL0 (hard coded)
    TXSYSCLKSEL                     => "00",   -- use PLL0 (hard coded)
    -- TX FPGA Interface Datapath Configuration
    TX8B10BEN                       => '1',
    -- GTPE2_CHANNEL Clocking
    PLL0CLK                         => pll0clk,
    PLL0REFCLK                      => pll0refclk,
    PLL1CLK                         => pll1clk,
    PLL1REFCLK                      => pll1refclk,
    -- Loopback
    LOOPBACK                        => loopback_i,
    -- PCI Express
    PHYSTATUS                       => open,
    RXRATE                          => "000",
    RXVALID                         => open,
    -- PMA Reserved
    PMARSVDIN3                      => '0',
    PMARSVDIN4                      => '0',
    -- Power-Down
    RXPD                            => powerdown_i,
    TXPD                            => powerdown_i,
    -- RX 8B/10B Decoder
    SETERRSTATUS                    => '0',
    -- RX Initialization and Reset
    EYESCANRESET                    => '0',
    RXUSERRDY                       => rxuserrdy_i,
    -- RX Margin Analysis
    EYESCANDATAERROR                => open,
    EYESCANMODE                     => '0',
    EYESCANTRIGGER                  => '0',
    -- RX Reset
    CLKRSVD0                        => '0',
    CLKRSVD1                        => '0',
    DMONFIFORESET                   => '0',
    DMONITORCLK                     => '0',
    RXPMARESETDONE                  => rxpmaresetdone,
    SIGVALIDCLK                     => '0',
    -- RX CDR
    RXCDRFREQRESET                  => '0',
    RXCDRHOLD                       => '0',
    RXCDRLOCK                       => open,
    RXCDROVRDEN                     => '0',
    RXCDRRESET                      => '0',
    RXCDRRESETRSV                   => '0',
    RXOSCALRESET                    => '0',
    RXOSINTCFG                      => "0010",
    RXOSINTDONE                     => open,
    RXOSINTHOLD                     => '0',
    RXOSINTOVRDEN                   => '0',
    RXOSINTPD                       => '0',
    RXOSINTSTARTED                  => open,
    RXOSINTSTROBE                   => '0',
    RXOSINTSTROBESTARTED            => open,
    RXOSINTTESTOVRDEN               => '0',
    --RX Clock Correction
    RXCLKCORCNT                     => open,
    -- RX FPGA Interface Datapath Configuration
    RX8B10BEN                       => '1',
    -- RX FPGA Interface
    RXDATA                          => rxdata,
    RXUSRCLK                        => usrclk,
    RXUSRCLK2                       => usrclk,
    -- RX Pattern Checker
    RXPRBSERR                       => open,
    RXPRBSSEL                       => "000",
    RXPRBSCNTRESET                  => '0',
    -- RX 8B/10B Decoder
    RXCHARISCOMMA                   => open,
    RXCHARISK                       => rxcharisk,
    RXDISPERR                       => rxdisperr,
    RXNOTINTABLE                    => rxnotintable,
    -- RX AFE
    GTPRXN                          => rxn_i,
    GTPRXP                          => rxp_i,
    PMARSVDIN2                      => '0',
    PMARSVDOUT0                     => open,
    PMARSVDOUT1                     => open,
    -- RX Buffer Bypass
    RXBUFRESET                      => '0',
    RXBUFSTATUS                     => rxbufstatus_o,
    RXDDIEN                         => '0',
    RXDLYBYPASS                     => '1',
    RXDLYEN                         => '0',
    RXDLYOVRDEN                     => '0',
    RXDLYSRESET                     => '0',
    RXDLYSRESETDONE                 => open,
    RXPHALIGN                       => '0',
    RXPHALIGNDONE                   => open,
    RXPHALIGNEN                     => '0',
    RXPHDLYPD                       => '0',
    RXPHDLYRESET                    => '0',
    RXPHMONITOR                     => open,
    RXPHOVRDEN                      => '0',
    RXPHSLIPMONITOR                 => open,
    RXSTATUS                        => open,
    RXSYNCALLIN                     => '0',
    RXSYNCDONE                      => open,
    RXSYNCIN                        => '0',
    RXSYNCMODE                      => '0',
    RXSYNCOUT                       => open,
    -- RX Byte and Word Alignment
    RXBYTEISALIGNED                 => rxbyteisaligned_o,
    RXBYTEREALIGN                   => rxbyterealign_o,
    RXCOMMADET                      => open, -- INFO: required for manual alignment
    RXCOMMADETEN                    => '1',  -- INFO: '0' for manual alignment
    RXMCOMMAALIGNEN                 => rxencommaalign_i,
    RXPCOMMAALIGNEN                 => rxencommaalign_i,
    RXSLIDE                         => '0',  -- INFO: required for manual alignment 
    -- RX Channel Bonding
    RXCHANBONDSEQ                   => open,
    RXCHBONDEN                      => '0',
    RXCHBONDI                       => "0000",
    RXCHBONDLEVEL                   => "000",
    RXCHBONDMASTER                  => '0',
    RXCHBONDO                       => open,
    RXCHBONDSLAVE                   => '0',
    -- RX Channel Bonding
    RXCHANISALIGNED                 => open,
    RXCHANREALIGN                   => open,
    -- RX Decision Feedback Equalizer (DFE)
    DMONITOROUT                     => open,
    RXADAPTSELTEST                  => "00000000000000",
    RXDFEXYDEN                      => '0',
    RXOSINTEN                       => '1',
    RXOSINTID0                      => "0000",
    RXOSINTNTRLEN                   => '0',
    RXOSINTSTROBEDONE               => open,
    -- RX Driver, OOB Signalling, Coupling and Equalizer, CDR
    RXLPMLFOVRDEN                   => '0',
    RXLPMOSINTNTRLEN                => '0',
    -- RX Equalizer
    RXLPMHFHOLD                     => '0',
    RXLPMHFOVRDEN                   => '0',
    RXLPMLFHOLD                     => '0',
    RXOSHOLD                        => '0',
    RXOSOVRDEN                      => '0',
    -- RX Fabric ClocK Output Control
    RXRATEDONE                      => open,
    RXRATEMODE                      => '0',
    RXOUTCLK                        => open,
    RXOUTCLKFABRIC                  => open,
    RXOUTCLKPCS                     => open,
    RXOUTCLKSEL                     => "010",
    -- RX Gearbox
    RXDATAVALID                     => open,
    RXHEADER                        => open,
    RXHEADERVALID                   => open,
    RXSTARTOFSEQ                    => open,
    RXGEARBOXSLIP                   => '0',
    -- RX Initialization and Reset
    GTRXRESET                       => rxreset,
    RXLPMRESET                      => '0',
    RXOOBRESET                      => '0',
    RXPCSRESET                      => '0',
    RXPMARESET                      => '0',
    -- RX OOB Signalling
    RXCOMSASDET                     => open,
    RXCOMWAKEDET                    => open,
    RXCOMINITDET                    => open,
    RXELECIDLE                      => open,
    RXELECIDLEMODE                  => "11",
    -- RX Polarity Control
    RXPOLARITY                      => '0',
    -- RX Initialization and Reset
    RXRESETDONE                     => rxresetdone_o,
    -- TX Buffer Bypass
    TXPHDLYTSTCLK                   => '0',
    -- TX Configurable Driver
    TXPOSTCURSOR                    => "00000",
    TXPOSTCURSORINV                 => '0',
    TXPRECURSOR                     => "00000",
    TXPRECURSORINV                  => '0',
    -- TX Fabric Clock Output Control
    TXRATEMODE                      => '0',
    -- TX Initialization and Reset
    CFGRESET                        => '0',
    GTTXRESET                       => txreset_i,
    PCSRSVDOUT                      => open,
    TXUSERRDY                       => txuserrdy_i,
    -- TX Phase Interpolator PPM Controller
    TXPIPPMEN                       => '0',
    TXPIPPMOVRDEN                   => '0',
    TXPIPPMPD                       => '0',
    TXPIPPMSEL                      => '1',
    TXPIPPMSTEPSIZE                 => "00000",
    -- Transceiver Reset Mode Operation
    GTRESETSEL                      => '0',
    RESETOVRD                       => '0',
    -- TX Reset
    TXPMARESETDONE                  => txpmaresetdone,
    -- TX Configurable Driver
    PMARSVDIN0                      => '0',
    PMARSVDIN1                      => '0',
    -- TX FPGA Interface
    TXDATA                          => txdata,
    TXUSRCLK                        => usrclk,
    TXUSRCLK2                       => usrclk,
    -- TX PCI Express
    TXELECIDLE                      => '0',
    TXMARGIN                        => "000",
    TXRATE                          => "000",
    TXSWING                         => '0',
    -- TX Pattern Generator
    TXPRBSFORCEERR                  => '0',
    -- TX 8B/10B Encoder
    TX8B10BBYPASS                   => "0000",
    TXCHARDISPMODE                  => "0000",
    TXCHARDISPVAL                   => "0000",
    TXCHARISK(3 downto 2)           => "00",
    TXCHARISK(1 downto 0)           => txcharisk_i,
    -- TX Buffer Bypass
    TXDLYBYPASS                     => '1',
    TXDLYEN                         => '0',
    TXDLYHOLD                       => '0',
    TXDLYOVRDEN                     => '0',
    TXDLYSRESET                     => '0',
    TXDLYSRESETDONE                 => open,
    TXDLYUPDOWN                     => '0',
    TXPHALIGN                       => '0',
    TXPHALIGNDONE                   => open,
    TXPHALIGNEN                     => '0',
    TXPHDLYPD                       => '0',
    TXPHDLYRESET                    => '0',
    TXPHINIT                        => '0',
    TXPHINITDONE                    => open,
    TXPHOVRDEN                      => '0',
    -- TX Buffer
    TXBUFSTATUS                     => open,
    -- TX Buffer and Phase Alignment
    TXSYNCALLIN                     => '0',
    TXSYNCDONE                      => open,
    TXSYNCIN                        => '0',
    TXSYNCMODE                      => '0',
    TXSYNCOUT                       => open,
    -- TX Configurable Driver
    GTPTXN                          => txn_o,
    GTPTXP                          => txp_o,
    TXBUFDIFFCTRL                   => "100",
    TXDEEMPH                        => '0',
    TXDIFFCTRL                      => "1000",
    TXDIFFPD                        => '0',
    TXINHIBIT                       => '0',
    TXMAINCURSOR                    => "0000000",
    TXPISOPD                        => '0',
    -- TX Fabric Clock Output Control
    TXOUTCLK                        => txoutclk,
    TXOUTCLKFABRIC                  => open,
    TXOUTCLKPCS                     => open,
    TXOUTCLKSEL                     => "010",
    TXRATEDONE                      => open,
    -- TX Gearbox
    TXGEARBOXREADY                  => open,
    TXHEADER                        => "000",
    TXSEQUENCE                      => "0000000",
    TXSTARTSEQ                      => '0',
    -- TX Initialization and Reset
    TXPCSRESET                      => '0',
    TXPMARESET                      => '0',
    TXRESETDONE                     => txresetdone_o,
    -- TX OOB Signalling
    TXCOMFINISH                     => open,
    TXCOMINIT                       => '0',
    TXCOMSAS                        => '0',
    TXCOMWAKE                       => '0',
    TXPDELECIDLEMODE                => '0',
    -- TX Polarity Control
    TXPOLARITY                      => '0',
    -- TX Receiver Detection
    TXDETECTRX                      => '0',
    -- TX Pattern Generator
    TXPRBSSEL                       => "000"
  );

  -- GTP reset sequence upon FPGA configuration (AR# 53561)
  -- Based on code generated by Vivado GT wizard (<gtname>_gtrxreset_seq.vhd)
  gen_gtrxreset_seq : if g_SIMULATION /= "TRUE" generate
    cmp_gtrxreset_seq_0 : gtrxreset_seq
    port map
    (
      RST             =>  init_rst_i,
      GTRXRESET_IN    =>  rxreset_i,
      RXPMARESETDONE  =>  rxpmaresetdone,
      GTRXRESET_OUT   =>  rxreset,
      DRP_OP_DONE     =>  drp_op_done,
      DRPCLK          =>  init_clk_i,
      DRPEN           =>  drpen,
      DRPADDR         =>  drpaddr,
      DRPWE           =>  drpwe,
      DRPDO           =>  drpdo,
      DRPDI           =>  drpdi,
      DRPRDY          =>  drprdy
    );
  end generate;

  gen_gtrxreset_seq_sim : if g_SIMULATION = "TRUE" generate
    cmp_gtrxreset_seq_0 : gtrxreset_seq_sim
    port map
    (
      RST             =>  init_rst_i,
      GTRXRESET_IN    =>  rxreset_i,
      RXPMARESETDONE  =>  rxpmaresetdone,
      GTRXRESET_OUT   =>  rxreset,
      DRP_OP_DONE     =>  drp_op_done,
      DRPCLK          =>  init_clk_i,
      DRPEN           =>  drpen,
      DRPADDR         =>  drpaddr,
      DRPWE           =>  drpwe,
      DRPDO           =>  drpdo,
      DRPDI           =>  drpdi,
      DRPRDY          =>  drprdy
    );
  end generate;

  -- Quad GTP PLL instance
  cmp_gtpll : GTPE2_COMMON
  generic map
  (
    -- Simulation
    SIM_RESET_SPEEDUP       => g_SIMULATION_SPEEDUP,
    SIM_PLL0REFCLK_SEL      => "001",
    SIM_PLL1REFCLK_SEL      => "001",
    SIM_VERSION             => "2.0",
    -- PLL Dividers
    PLL0_FBDIV              => c_PLLFBDIV,
    PLL0_FBDIV_45           => c_PLLFBDIV45,
    PLL0_REFCLK_DIV         => c_PLLREFDIV,
    PLL1_FBDIV              => 1,
    PLL1_FBDIV_45           => 4,
    PLL1_REFCLK_DIV         => 1,
    -- Common Block
    BIAS_CFG                => x"0000000000050001",
    COMMON_CFG              => x"00000000",
    -- PLL
    PLL0_CFG                => x"01F03DC",
    PLL0_DMON_CFG           => '0',
    PLL0_INIT_CFG           => x"00001E",
    PLL0_LOCK_CFG           => x"1E8",
    PLL1_CFG                => x"01F03DC",
    PLL1_DMON_CFG           => '0',
    PLL1_INIT_CFG           => x"00001E",
    PLL1_LOCK_CFG           => x"1E8",
    PLL_CLKOUT_CFG          => x"00",
    -- Reserved
    RSVD_ATTR0              => x"0000",
    RSVD_ATTR1              => x"0000"
  )
  port map
  (
    DMONITOROUT             => open,
    -- Dynamic Reconfiguration Port (DRP)
    DRPADDR                 => "00000000",
    DRPCLK                  => '0',
    DRPDI                   => "0000000000000000",
    DRPDO                   => open,
    DRPEN                   => '0',
    DRPRDY                  => open,
    DRPWE                   => '0',
    -- GTPE2_COMMON Clocking
    GTGREFCLK0              => '0',
    GTGREFCLK1              => '0',
    GTEASTREFCLK0           => '0',
    GTEASTREFCLK1           => '0',
    GTREFCLK0               => refclk0_i,
    GTREFCLK1               => refclk1_i,
    GTWESTREFCLK0           => '0',
    GTWESTREFCLK1           => '0',
    PLL0OUTCLK              => pll0clk,
    PLL0OUTREFCLK           => pll0refclk,
    PLL1OUTCLK              => pll1clk,
    PLL1OUTREFCLK           => pll1refclk,
    -- PLL                  
    PLL0FBCLKLOST           => open,
    PLL0LOCK                => pll_lock_o,
    PLL0LOCKDETCLK          => pll_lockdetclk_i,
    PLL0LOCKEN              => '1',
    PLL0PD                  => '0',
    PLL0REFCLKLOST          => pll_refclklost_o,
    PLL0REFCLKSEL           => pll_refclksel_i,
    PLL0RESET               => pll_rst_i,
    PLL1FBCLKLOST           => open,
    PLL1LOCK                => open,
    PLL1LOCKDETCLK          => '0',
    PLL1LOCKEN              => '1',
    PLL1PD                  => '1',
    PLL1REFCLKLOST          => open,
    PLL1REFCLKSEL           => "001",
    PLL1RESET               => '0',
    -- Common Block         
    BGRCALOVRDENB           => '1',
    PLLRSVD1                => "0000000000000000",
    PLLRSVD2                => "00000",
    REFCLKOUTMONITOR0       => open,
    REFCLKOUTMONITOR1       => open,
    -- RX AFE               
    PMARSVDOUT              => open,
    -- QPLL                 
    BGBYPASSB               => '1',
    BGMONITORENB            => '1',
    BGPDB                   => '1',
    BGRCALOVRD              => "11111",
    PMARSVD                 => "00000000",
    RCALENB                 => '1'
  );

  -- User clock global buffer
  txoutclk_bufg0_i : BUFG
  port map
  (
    I       => txoutclk,
    O       => usrclk
  );

  usrclk_o <= usrclk;

end rtl;
