//-----------------------------------------------------------------------------
// Title      : GTPE2 RX elastic buffer testbench
// Project    : Open Communication Controller
//-----------------------------------------------------------------------------
// Author     : Daniel Tavares
// Company    : CNPEM LNLS-DIG
// Created    : 2020-05-08
// Platform   : Xilinx
//-----------------------------------------------------------------------------
// Copyright (c) 2020 CNPEM
//
// This source describes open hardware and is licensed under the CERN-OHL-W v2.
//
// You may redistribute and modify this documentation and make products using
// it under the terms of the CERN-OHL-W v2 (https:/cern.ch/cern-ohl), or (at
// your option) any later version. This documentation is distributed WITHOUT
// ANY EXPRESS OR IMPLIED WARRANTY, INCLUDING OF MERCHANTABILITY, SATISFACTORY
// QUALITY AND FITNESS FOR A PARTICULAR PURPOSE. Please see the CERN-OHL-W v2
// for applicable conditions.
//-----------------------------------------------------------------------------

`timescale 1ns / 1ps

module main;

  //------------
  // Parameters
  //------------
  localparam REFCLK_PERIOD = 8.0;               // [ns]
  localparam USRCLK_PERIOD = REFCLK_PERIOD/2.5; // [ns]
  localparam INITCLK_PERIOD = 10.0;             // [ns]
  localparam BLIND_PERIOD = 10;                 // [usrclk cycles]
  localparam PLLRST_PERIOD = 2500;              // [refclk cycles]
  localparam IDLE_PERIOD = 193;                 // [usrclk cycles]
  localparam NUM_TRIES = 10;
  localparam NUM_SUCCESFUL_DATA = 1000;
  localparam IDLE = 16'hbc95;

  //---------
  // Signals
  //---------
  reg refclk = 0;
  reg pll_rst = 0;
  reg rxreset = 0;
  reg txreset = 0;
  reg rxuserrdy = 1;
  reg txuserrdy = 1;
  wire rxencommaalign;
  wire [1:0]  txcharisk;
  wire [15:0] txdata;
  reg pll_lock_reg;
  wire usrclk;
  wire rxtxn, rxtxp;
  wire rxbyteisaligned;
  wire [1:0] rxcharisk, rxdisperr, rxnotintable;
  wire [2:0] rxbufstatus;
  wire [15:0] rxdata;
  wire rxresetdone;
  wire txresetdone;
  wire pll_lock;
  reg rdy;
  wire fail;
  
  wire [31:0] latency_min;
  wire [31:0] latency_max;
  integer cnt_tries;
  
  //--------
  // Clocks
  //--------
  always begin
    refclk = ~refclk;
    #(REFCLK_PERIOD/2);
  end

  //-------------------------------
  // Resets and Simulation control
  //------------------------------
  initial begin
    // Keep reseting the whole design by NUM_TRIES times
    for (cnt_tries = 1; cnt_tries <= NUM_TRIES; cnt_tries = cnt_tries + 1) begin
      $display("Reset try #%.3d...", cnt_tries);

      pll_rst = 1;
      #(200*REFCLK_PERIOD);
      pll_rst = 0;
      #((PLLRST_PERIOD-200)*REFCLK_PERIOD);

      if (!fail) begin
        $display("Latency [txuserclk cycles]: %d (min) - %d (max).", latency_min, latency_max);
        $display("PASS");
        $finish;
      end
    end
    $display("FAIL");
    $finish;
  end

  //--------------------
  // GTP reset sequence
  //--------------------
  always @(posedge refclk) begin
    // Pulse GTP reset and set RX and TX user ready signals once GTP PLL lock
    // has been achieved. Note this must be done in refclk domain, not usrclk
    // domain since usrclk is generated by the GTP itself, thus unavailable
    // during reset.
    pll_lock_reg <= pll_lock;
    rxreset <= pll_lock ^ pll_lock_reg;
    txreset <= pll_lock ^ pll_lock_reg;

    if (pll_lock == 1) begin
      rxuserrdy <= 1;
      txuserrdy <= 1;
    end  
    else if (pll_lock == 0) begin
      rxuserrdy <= 0;
      txuserrdy <= 0;
    end

    rdy <= rxuserrdy && txuserrdy && rxresetdone && txresetdone;
  end

  //-------------------
  // Design validation
  //-------------------
  rxbuffer_checker #
  (
    .g_IDLE                 (IDLE),
    .g_IDLE_PERIOD          (IDLE_PERIOD),
    .g_NUM_TRIES            (NUM_TRIES),
    .g_BLIND_PERIOD         (BLIND_PERIOD),
    .g_NUM_SUCCESFUL_DATA   (NUM_SUCCESFUL_DATA)
  )
  cmp_latency_checker
  (
    .fail_o             (fail),
    .usrclk_i           (usrclk),
    .valid_i            (rdy),
    .rx_data_i          (rxdata),
    .rx_k_i             (rxcharisk),
    .tx_data_i          (txdata),
    .tx_k_i             (txcharisk),
    .rx_realign_o       (rxencommaalign),
    .rx_aligned_o       (rxbyteisaligned),
    .rx_bufstatus_i     (rxbufstatus),
    .latency_min_o      (latency_min),
    .latency_max_o      (latency_max)
  );

  // ----
  // DUT 
  // ----
  occ_gtpe2_tile #(
    .g_SIMULATION           ("TRUE"),
    .g_SIMULATION_SPEEDUP   ("TRUE")
  )
  cmp_occ_gtpe2_tile (
    .rxn_i              (rxtxn),
    .rxp_i              (rxtxp),
    .txn_o              (rxtxn),
    .txp_o              (rxtxp),
    .rxreset_i          (rxreset),
    .rxresetdone_o      (rxresetdone),
    .rxcharisk_o        (rxcharisk),
    .rxdisperr_o        (rxdisperr),
    .rxnotintable_o     (rxnotintable),
    .rxbyteisaligned_o  (rxbyteisaligned),
    .rxbyterealign_o    (rxbyterealign),
    .rxencommaalign_i   (rxencommaalign),
    .rxbufstatus_o      (rxbufstatus),
    .rxdata_o           (rxdata),
    .rxuserrdy_i        (rxuserrdy),
    .txreset_i          (txreset),
    .txresetdone_o      (txresetdone),
    .txcharisk_i        (txcharisk),
    .txdata_i           (txdata),
    .txuserrdy_i        (txuserrdy),
    .refclk0_i          (refclk),
    .refclk1_i          (refclk),
    .usrclk_o           (usrclk),
    .loopback_i         (3'b000),
    .powerdown_i        (2'b00),
    .pll_lockdetclk_i   (refclk),
    .pll_lock_o         (pll_lock),
    .pll_refclklost_o   (),
    .pll_refclksel_i    (3'b001),
    .pll_rst_i          (pll_rst),
    .init_rst_i         (1'b0),
    .init_clk_i         (refclk)
  );

endmodule
