//-----------------------------------------------------------------------------
// Title      : GTPE2 RX elastic buffer testbench
// Project    : Open Communication Controller
//-----------------------------------------------------------------------------
// Author     : Daniel Tavares
// Company    : CNPEM LNLS-DIG
// Created    : 2020-05-08
// Platform   : Xilinx
//-----------------------------------------------------------------------------
// Copyright (c) 2020 CNPEM
//
// This source describes open hardware and is licensed under the CERN-OHL-W v2.
//
// You may redistribute and modify this documentation and make products using
// it under the terms of the CERN-OHL-W v2 (https:/cern.ch/cern-ohl), or (at
// your option) any later version. This documentation is distributed WITHOUT
// ANY EXPRESS OR IMPLIED WARRANTY, INCLUDING OF MERCHANTABILITY, SATISFACTORY
// QUALITY AND FITNESS FOR A PARTICULAR PURPOSE. Please see the CERN-OHL-W v2
// for applicable conditions.
//-----------------------------------------------------------------------------

`timescale 1ns / 1ps

module main;

  //------------
  // Parameters
  //------------
  localparam REFCLK_PERIOD = 8.0;               // [ns]
  localparam USRCLK_PERIOD = REFCLK_PERIOD/2.5; // [ns]
  localparam INITCLK_PERIOD = 10.0;             // [ns]
  localparam BLIND_PERIOD = 10;                 // [usrclk cycles]
  localparam PLLRST_PERIOD = 2500;              // [refclk cycles]
  localparam IDLE_PERIOD = 193;                 // [usrclk cycles]
  localparam NUM_TRIES = 10;
  localparam NUM_SUCCESFUL_DATA = 1000;
  localparam IDLE = 16'hbc95;

  //---------
  // Signals
  //---------
  reg refclk = 0;
  reg pll_rst = 0;
  reg rxreset = 0;
  reg txreset = 0;
  reg rxuserrdy = 1;
  reg txuserrdy = 1;
  reg rxencommaalign;
  reg [1:0]  txcharisk;
  reg [15:0] txdata;
  reg pll_lock_reg;
  reg right_comma_byte = 0;
  wire usrclk;
  wire rxtxn, rxtxp;
  wire rxbyteisaligned;
  wire [1:0] rxcharisk, rxdisperr, rxnotintable;
  wire [2:0] rxbufstatus;
  wire [15:0] rxdata;
  wire rxresetdone;
  wire txresetdone;
  wire pll_lock;

  integer latency = 0;
  integer latency_min = 100000;
  integer latency_max = 0;

  integer cnt_data = 0;
  integer cnt_blind = 0;
  integer cnt_tries = 1;
  integer cnt_succesful_data = 0;
  
  //--------
  // Clocks
  //--------
  always begin
    refclk = ~refclk;
    #(REFCLK_PERIOD/2);
  end

  //--------
  // Resets
  //--------
  initial begin
    // Keep reseting the whole system and tracking number of tries
    forever begin
      pll_rst = 1;
      #(200*REFCLK_PERIOD);
      pll_rst = 0;
      #((PLLRST_PERIOD-200)*REFCLK_PERIOD);
      cnt_tries = cnt_tries + 1;
    end
  end

  //--------------------
  // GTP reset sequence
  //--------------------
  always @(posedge refclk) begin
    // Pulse GTP reset and set RX and TX user ready signals once GTP PLL lock
    // has been achieved. Note this must be done in refclk domain, not usrclk
    // domain since usrclk is generated by the GTP itself, thus unavailable
    // during reset.
    pll_lock_reg <= pll_lock;
    rxreset <= pll_lock ^ pll_lock_reg;
    txreset <= pll_lock ^ pll_lock_reg;

    if (pll_lock == 1) begin
      rxuserrdy <= 1;
      txuserrdy <= 1;
    end  
    else if (pll_lock == 0) begin
      rxuserrdy <= 0;
      txuserrdy <= 0;
    end
  end

  //-----------------
  // Data generation
  //-----------------
  always @(posedge usrclk) begin
    // Produce data incremented by 1 in order to allow latency calculation
    // Interleave with IDLE words for comma alignment and clock correction
    if (cnt_data % IDLE_PERIOD == 0) begin
      txcharisk <= 2'b10;
      txdata <= IDLE;
    end
    else begin
      txcharisk <= 2'b00;
      txdata <= cnt_data;
    end
    cnt_data = cnt_data + 1;
  end

  //-------------------
  // Design validation
  //-------------------
  always @(posedge usrclk) begin
    if (rxuserrdy == 1 && txuserrdy == 1 && rxresetdone == 1 && txresetdone == 1) begin
      rxencommaalign <= 1;
    end
    else if (rxuserrdy == 0 || txuserrdy == 0 || rxbyteisaligned == 1) begin
      rxencommaalign <= 0;
    end

    if (rxbyteisaligned == 1) begin
      if (cnt_blind > BLIND_PERIOD) begin
        // The blind period is used to ignore the first cycles after the GTP
        // signals that the comma alignment has been achieved through the
        // rxbyteisaligned port. UG482 is not clear about how many clock cycles
        // it takes for data coming out at the rxdata port is guaranteed to be
        // aligned as indicated by rxbyteisaligned.
        if (rxcharisk == 2'b00) begin
          if (right_comma_byte == 1) begin
            // Data is byte-aligned - Receiveing payload
            if (txcharisk == 2'b00) begin
              // When TX and RX data have no K character it is possible to
              // calculate overall TX-RX latency - it must be assured the comma
              // byte alignment have been already performed
              latency = txdata - rxdata;
              cnt_succesful_data = cnt_succesful_data + 1;

              // Latency statistics
              if (latency > latency_max) latency_max = latency;
              if (latency < latency_min) latency_min = latency;        

              if (cnt_succesful_data > NUM_SUCCESFUL_DATA) begin
                $display("Latency [txuserclk cycles]: %d (min) - %d (max).", latency_min, latency_max);
                $display("PASS");
                $finish;
              end
            end
          end
        end
        else if (rxcharisk == 2'b10 && rxdata == IDLE) begin
          // Data is byte-aligned - Comma in the right byte of an IDLE word
          right_comma_byte = 1;
        end
        else if (rxcharisk == 2'b01 && rxdata[7:0] == IDLE[15:8]) begin
          // Data is not byte-aligned - Comma in the wrong byte of an IDLE word
            if (cnt_tries >= NUM_TRIES) begin
              $display("Wrong comma byte alignment. Number of reset tries: %d.", NUM_TRIES);
              $display("FAIL");
              $stop;
            end
        end
        else begin
          if (cnt_tries >= NUM_TRIES) begin
            $display("Unknown comma misalignment. Number of reset tries: %d.", NUM_TRIES);
            $display("FAIL");
            $stop;
          end
        end
      end
      cnt_blind = cnt_blind + 1;
    end
    else begin
      cnt_blind = 0;
      right_comma_byte = 0;
    end
  end

  // ----
  // DUT 
  // ----
  occ_gtpe2_tile #(
    .g_SIMULATION           ("TRUE"),
    .g_SIMULATION_SPEEDUP   ("TRUE")
  )
  cmp_occ_gtpe2_tile (
    .rxn_i              (rxtxn),
    .rxp_i              (rxtxp),
    .txn_o              (rxtxn),
    .txp_o              (rxtxp),
    .rxreset_i          (rxreset),
    .rxresetdone_o      (rxresetdone),
    .rxcharisk_o        (rxcharisk),
    .rxdisperr_o        (rxdisperr),
    .rxnotintable_o     (rxnotintable),
    .rxbyteisaligned_o  (rxbyteisaligned),
    .rxbyterealign_o    (rxbyterealign),
    .rxencommaalign_i   (rxencommaalign),
    .rxbufstatus_o      (rxbufstatus),
    .rxdata_o           (rxdata),
    .rxuserrdy_i        (rxuserrdy),
    .txreset_i          (txreset),
    .txresetdone_o      (txresetdone),
    .txcharisk_i        (txcharisk),
    .txdata_i           (txdata),
    .txuserrdy_i        (txuserrdy),
    .refclk0_i          (refclk),
    .refclk1_i          (refclk),
    .usrclk_o           (usrclk),
    .loopback_i         (3'b000),
    .powerdown_i        (2'b00),
    .pll_lockdetclk_i   (refclk),
    .pll_lock_o         (pll_lock),
    .pll_refclklost_o   (),
    .pll_refclksel_i    (3'b001),
    .pll_rst_i          (pll_rst),
    .init_rst_i         (1'b0),
    .init_clk_i         (refclk)
  );

endmodule
