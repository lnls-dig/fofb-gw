-------------------------------------------------------------------------------
-- Title      : Xilinx 7-series GTP Transceiver with OCC configurations
-- Project    : Open Communication Controller
-------------------------------------------------------------------------------
-- Author     : Daniel Tavares
-- Company    : CNPEM LNLS-DIG
-- Created    : 2020-05-18
-- Platform   : Xilinx
-------------------------------------------------------------------------------
-- Description: Encapsulates Xilinx 7-series GTP transceiver and corresponding
-- PLL and clock buffers with the settings required by the Open Communication
-- Controller protocol. One tile instance comprehends 1 to 4 transceivers.
--
-- Based on code generated by Vivado GT wizard (gtrxreset_seq.vhd) for the
-- receiver reset sequence (AR# 53561).
-------------------------------------------------------------------------------
--
-- Copyright (c) 2020 CNPEM
--
-- This source describes open hardware and is licensed under the CERN-OHL-W v2.
--
-- You may redistribute and modify this documentation and make products using
-- it under the terms of the CERN-OHL-W v2 (https:/cern.ch/cern-ohl, or (at
-- your option) any later version. This documentation is distributed WITHOUT
-- ANY EXPRESS OR IMPLIED WARRANTY, INCLUDING OF MERCHANTABILITY, SATISFACTORY
-- QUALITY AND FITNESS FOR A PARTICULAR PURPOSE. Please see the CERN-OHL-W v2
-- for applicable conditions.
--
-------------------------------------------------------------------------------

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

-- Synchronizers
use work.gencores_pkg.all;

library unisim;
use unisim.vcomponents.all;

entity occ_gtp_phy_family7 is
generic
(
  g_SIMULATION        : string               := "FALSE";
  g_NUM_CHANNELS      : integer range 1 to 4 := 1;          -- TODO: g_NUM_CHANNELS should range from 1 to 4
  g_REFCLK            : string               := "REFCLK0"   -- TODO: select among "REFCLK0", "REFCLK1", "EASTREFCLK0", "EASTREFCLK1", "WESTREFCLK0", "WESTREFCLK1"
);
port
(
  -----------------
  -- EXTERNAL PADS
  -----------------
  pad_txn_o       : out std_logic;
  pad_txp_o       : out std_logic;
  pad_rxn_i       : in  std_logic;
  pad_rxp_i       : in  std_logic;
  pad_refclkn_i   : in  std_logic;
  pad_refclkp_i   : in  std_logic;

  ------------------
  -- INITIALIZATION
  ------------------
  rst_i           : in  std_logic;

  --------------------
  -- TRANSMITTER (TX)
  --------------------
  tx_rst_i        : in  std_logic;
  tx_clk_o        : out std_logic;
  tx_data_i       : in  std_logic_vector(15 downto 0);
  tx_k_i          : in  std_logic_vector(1 downto 0);
  tx_rdy_o        : out std_logic;

  -----------------
  -- RECEIVER (RX)
  -----------------
  rx_rst_i        : in  std_logic;
  rx_clk_o        : out std_logic;
  rx_data_o       : out std_logic_vector(15 downto 0);
  rx_k_o          : out std_logic_vector(1 downto 0);
  rx_resync_i     : in  std_logic;
  rx_synced_o     : out std_logic;
  rx_rdy_o        : out std_logic;
  rx_enc_err_o    : out std_logic;
  rx_buf_err_o    : out std_logic;

  -----------------
  -- CONFIGURATION
  -----------------
  loopen_i        : in  std_logic_vector(2 downto 0)
);
end occ_gtp_phy_family7;

architecture rtl of occ_gtp_phy_family7 is
  -- Reset wait time in number of refclk cycles (must be greater than 500 ns)
  constant c_RST_DELAY        : integer := 300;

  -- PLL dividers configuration
  constant c_PLLFBDIV         : integer := 5;
  constant c_PLLFBDIV45       : integer := 5;
  constant c_PLLREFDIV        : integer := 1;

  -- PLL reset and clock signals
  signal pll_lock             : std_logic;
  signal pll_rst              : std_logic;
  signal ref_clk              : std_logic;

  signal gteastrefclk0        : std_logic;
  signal gteastrefclk1        : std_logic;
  signal gtrefclk0            : std_logic;
  signal gtrefclk1            : std_logic;
  signal gtwestrefclk0        : std_logic;
  signal gtwestrefclk1        : std_logic;

  signal pll0refclksel        : std_logic_vector(2 downto 0);
  signal pll0clk              : std_logic;
  signal pll0refclk           : std_logic;
  signal pll1clk              : std_logic;
  signal pll1refclk           : std_logic;  

  -- Reset-related signals
  signal rst_synced           : std_logic;

  signal rx_rst               : std_logic;
  signal rx_rst_done          : std_logic;

  signal tx_rst               : std_logic;
  signal tx_rst_done          : std_logic;

  -- RX datapath signals
  signal rx_data_full         : std_logic_vector(31 downto 0);
  signal rx_k_full            : std_logic_vector(3 downto 0);
  signal rx_disp_err          : std_logic_vector(3 downto 0);
  signal rx_code_err          : std_logic_vector(3 downto 0);
  signal rx_clk               : std_logic;

  -- TX datapath signals and clocks
  signal tx_data_full         : std_logic_vector(31 downto 0);
  signal tx_clk_bufin         : std_logic;
  signal tx_clk               : std_logic;

  -- RX Elastic Buffer
  signal rx_bufstatus         : std_logic_vector(2 downto 0);

  -- RX reset sequence signals (AR# 53561)
  signal rx_pma_rst_done      : std_logic;
  signal tx_pma_rst_done      : std_logic;
  signal rx_rst_seqout        : std_logic;
  signal drp_done             : std_logic;
  signal drp_addr             : std_logic_vector(8 downto 0);
  signal drp_en               : std_logic;
  signal drp_we               : std_logic;
  signal drp_dataout          : std_logic_vector(15 downto 0);
  signal drp_datain           : std_logic_vector(15 downto 0);
  signal drp_rdy              : std_logic;

  -- RX reset sequence component (AR# 53561)
  component gtrxreset_seq_sim
  port ( 
    RST             : in  std_logic;
    GTRXRESET_IN    : in  std_logic;
    RXPMARESETDONE  : in  std_logic;
    GTRXRESET_OUT   : out std_logic;  
    DRPCLK          : in  std_logic;
    DRPADDR         : out std_logic_vector(8 downto 0);
    DRPDO           : in  std_logic_vector(15 downto 0);
    DRPDI           : out std_logic_vector(15 downto 0);
    DRPRDY          : in  std_logic;
    DRPEN           : out std_logic;
    DRPWE           : out std_logic;
    DRP_OP_DONE     : out std_logic
  );
  end component;

  component gtrxreset_seq
  port ( 
    RST             : in  std_logic;
    GTRXRESET_IN    : in  std_logic;
    RXPMARESETDONE  : in  std_logic;
    GTRXRESET_OUT   : out std_logic;  
    DRPCLK          : in  std_logic;
    DRPADDR         : out std_logic_vector(8 downto 0);
    DRPDO           : in  std_logic_vector(15 downto 0);
    DRPDI           : out std_logic_vector(15 downto 0);
    DRPRDY          : in  std_logic;
    DRPEN           : out std_logic;
    DRPWE           : out std_logic;
    DRP_OP_DONE     : out std_logic
  );
  end component;

begin

  -- GTPE2_CHANNEL instances
  cmp_gtpe2_0 : GTPE2_CHANNEL
  generic map
  (
    -- Simulation
    SIM_RECEIVER_DETECT_PASS        => "TRUE",
    SIM_RESET_SPEEDUP               => g_SIMULATION,
    SIM_TX_EIDLE_DRIVE_LEVEL        => "X",
    SIM_VERSION                     => "2.0",
    -- RX Byte and Word Alignment   
    ALIGN_COMMA_DOUBLE              => "FALSE",
    ALIGN_COMMA_ENABLE              => "1111111111",
    ALIGN_COMMA_WORD                => 2,
    ALIGN_MCOMMA_DET                => "TRUE",
    ALIGN_MCOMMA_VALUE              => "1010000011", -- -K28.5+ (10-bit symbol)
    ALIGN_PCOMMA_DET                => "TRUE",
    ALIGN_PCOMMA_VALUE              => "0101111100", -- +K28.5- (10-bit symbol)
    SHOW_REALIGN_COMMA              => "FALSE",
    RXSLIDE_AUTO_WAIT               => 7,
    RXSLIDE_MODE                    => "OFF",
    RX_SIG_VALID_DLY                => 10,
    -- RX 8B/10B Decoder            
    RX_DISPERR_SEQ_MATCH            => "TRUE",
    DEC_MCOMMA_DETECT               => "TRUE",
    DEC_PCOMMA_DETECT               => "TRUE",
    DEC_VALID_COMMA_ONLY            => "FALSE",
    -- RX Clock Correction          
    CBCC_DATA_SOURCE_SEL            => "DECODED",
    CLK_COR_SEQ_2_USE               => "FALSE",
    CLK_COR_KEEP_IDLE               => "FALSE",
    CLK_COR_MAX_LAT                 => 15,
    CLK_COR_MIN_LAT                 => 12,
    CLK_COR_PRECEDENCE              => "TRUE",
    CLK_COR_REPEAT_WAIT             => 0,
    CLK_COR_SEQ_LEN                 => 2,
    CLK_COR_SEQ_1_ENABLE            => "1111",
    CLK_COR_SEQ_1_1                 => "0110111100", -- K28.5 (8-bit symbol)
    CLK_COR_SEQ_1_2                 => "0010010101", -- D21.4 (8-bit symbol)
    CLK_COR_SEQ_1_3                 => "0000000000",
    CLK_COR_SEQ_1_4                 => "0000000000",
    CLK_CORRECT_USE                 => "TRUE",
    CLK_COR_SEQ_2_ENABLE            => "1111",
    CLK_COR_SEQ_2_1                 => "0000000000",
    CLK_COR_SEQ_2_2                 => "0000000000",
    CLK_COR_SEQ_2_3                 => "0000000000",
    CLK_COR_SEQ_2_4                 => "0000000000",
    -- RX Channel Bonding           
    CHAN_BOND_KEEP_ALIGN            => "FALSE",
    CHAN_BOND_MAX_SKEW              => 1,
    CHAN_BOND_SEQ_LEN               => 1,
    CHAN_BOND_SEQ_1_1               => "0000000000",
    CHAN_BOND_SEQ_1_2               => "0000000000",
    CHAN_BOND_SEQ_1_3               => "0000000000",
    CHAN_BOND_SEQ_1_4               => "0000000000",
    CHAN_BOND_SEQ_1_ENABLE          => "1111",
    CHAN_BOND_SEQ_2_1               => "0000000000",
    CHAN_BOND_SEQ_2_2               => "0000000000",
    CHAN_BOND_SEQ_2_3               => "0000000000",
    CHAN_BOND_SEQ_2_4               => "0000000000",
    CHAN_BOND_SEQ_2_ENABLE          => "1111",
    CHAN_BOND_SEQ_2_USE             => "FALSE",
    FTS_DESKEW_SEQ_ENABLE           => "1111",
    FTS_LANE_DESKEW_CFG             => "1111",
    FTS_LANE_DESKEW_EN              => "FALSE",
    -- RX Margin Analysis           
    ES_CONTROL                      => "000000",
    ES_ERRDET_EN                    => "FALSE",
    ES_EYE_SCAN_EN                  => "FALSE",
    ES_HORZ_OFFSET                  => x"010",
    ES_PMA_CFG                      => "0000000000",
    ES_PRESCALE                     => "00000",
    ES_QUALIFIER                    => x"00000000000000000000",
    ES_QUAL_MASK                    => x"00000000000000000000",
    ES_SDATA_MASK                   => x"00000000000000000000",
    ES_VERT_OFFSET                  => "000000000",
    -- RX FPGA Interface            
    RX_DATA_WIDTH                   => 20,
    -- PMA                          
    OUTREFCLK_SEL_INV               => "11",
    PMA_RSV                         => x"00000333",
    PMA_RSV2                        => x"00002040",
    PMA_RSV3                        => "00",
    PMA_RSV4                        => "0000",
    RX_BIAS_CFG                     => "0000111100110011",
    DMONITOR_CFG                    => x"000A00",
    RX_CM_SEL                       => "01",
    RX_CM_TRIM                      => "0000",
    RX_DEBUG_CFG                    => "00000000000000",
    RX_OS_CFG                       => "0000010000000",
    TERM_RCAL_CFG                   => "100001000010000",
    TERM_RCAL_OVRD                  => "000",
    TST_RSV                         => x"00000000",
    RX_CLK25_DIV                    => 5, -- TODO: operates for refclk up to 125 MHz only? Look at UG196
    TX_CLK25_DIV                    => 5, -- TODO: operates for refclk up to 125 MHz only? Look at UG196
    UCODEER_CLR                     => '0',
    -- PCI Express                  
    PCS_PCIE_EN                     => "FALSE",
    -- PCS                          
    PCS_RSVD_ATTR                   => x"000000000000",
    -- RX Buffer                    
    RXBUF_ADDR_MODE                 => "FULL",
    RXBUF_EIDLE_HI_CNT              => "1000",
    RXBUF_EIDLE_LO_CNT              => "0000",
    RXBUF_EN                        => "TRUE",
    RX_BUFFER_CFG                   => "000000",
    RXBUF_RESET_ON_CB_CHANGE        => "TRUE",
    RXBUF_RESET_ON_COMMAALIGN       => "FALSE",
    RXBUF_RESET_ON_EIDLE            => "FALSE",
    RXBUF_RESET_ON_RATE_CHANGE      => "TRUE",
    RXBUFRESET_TIME                 => "00001",
    RXBUF_THRESH_OVFLW              => 61,
    RXBUF_THRESH_OVRD               => "FALSE",
    RXBUF_THRESH_UNDFLW             => 4,
    RXDLY_CFG                       => x"001F",
    RXDLY_LCFG                      => x"030",
    RXDLY_TAP_CFG                   => x"0000",
    RXPH_CFG                        => x"C00002",
    RXPHDLY_CFG                     => x"084020",
    RXPH_MONITOR_SEL                => "00000",
    RX_XCLK_SEL                     => "RXREC",
    RX_DDI_SEL                      => "000000",
    RX_DEFER_RESET_BUF_EN           => "TRUE",
    -- CDR                          
    RXCDR_CFG                       => x"0000107FE406001041010", -- INFO: depends on RXOUT_DIV attribute
    RXCDR_FR_RESET_ON_EIDLE         => '0',
    RXCDR_HOLD_DURING_EIDLE         => '0',
    RXCDR_PH_RESET_ON_EIDLE         => '0',
    RXCDR_LOCK_CFG                  => "001001",
    -- RX Initialization and Reset  
    RXCDRFREQRESET_TIME             => "00001",
    RXCDRPHRESET_TIME               => "00001",
    RXISCANRESET_TIME               => "00001",
    RXPCSRESET_TIME                 => "00001",
    RXPMARESET_TIME                 => "00011",
    -- RX OOB Signalling            
    RXOOB_CFG                       => "0000110",
    -- RX Gearbox                   
    RXGEARBOX_EN                    => "FALSE",
    GEARBOX_MODE                    => "000",
    -- PRBS Detection               
    RXPRBS_ERR_LOOPBACK             => '0',
    -- Power-Down                   
    PD_TRANS_TIME_FROM_P2           => x"03c",
    PD_TRANS_TIME_NONE_P2           => x"3c",
    PD_TRANS_TIME_TO_P2             => x"64",
    -- RX OOB Signalling            
    SAS_MAX_COM                     => 64,
    SAS_MIN_COM                     => 36,
    SATA_BURST_SEQ_LEN              => "0101",
    SATA_BURST_VAL                  => "100",
    SATA_EIDLE_VAL                  => "100",
    SATA_MAX_BURST                  => 8,
    SATA_MAX_INIT                   => 21,
    SATA_MAX_WAKE                   => 7,
    SATA_MIN_BURST                  => 4,
    SATA_MIN_INIT                   => 12,
    SATA_MIN_WAKE                   => 4,
    -- RX Fabric Clock Output Control
    TRANS_TIME_RATE                 => x"0E",
    -- TX Buffer                    
    TXBUF_EN                        => "TRUE",
    TXBUF_RESET_ON_RATE_CHANGE      => "TRUE",
    TXDLY_CFG                       => x"001F",
    TXDLY_LCFG                      => x"030",
    TXDLY_TAP_CFG                   => x"0000",
    TXPH_CFG                        => x"0780",
    TXPHDLY_CFG                     => x"084020",
    TXPH_MONITOR_SEL                => "00000",
    TX_XCLK_SEL                     => "TXOUT",
    -- TX FPGA Interface            
    TX_DATA_WIDTH                   => 20,
    -- TX Configurable Driver       
    TX_DEEMPH0                      => "000000",
    TX_DEEMPH1                      => "000000",
    TX_EIDLE_ASSERT_DELAY           => "110",
    TX_EIDLE_DEASSERT_DELAY         => "100",
    TX_LOOPBACK_DRIVE_HIZ           => "FALSE",
    TX_MAINCURSOR_SEL               => '0',
    TX_DRIVE_MODE                   => "DIRECT",
    TX_MARGIN_FULL_0                => "1001110",
    TX_MARGIN_FULL_1                => "1001001",
    TX_MARGIN_FULL_2                => "1000101",
    TX_MARGIN_FULL_3                => "1000010",
    TX_MARGIN_FULL_4                => "1000000",
    TX_MARGIN_LOW_0                 => "1000110",
    TX_MARGIN_LOW_1                 => "1000100",
    TX_MARGIN_LOW_2                 => "1000010",
    TX_MARGIN_LOW_3                 => "1000000",
    TX_MARGIN_LOW_4                 => "1000000",
    -- TX Gearbox                   
    TXGEARBOX_EN                    => "FALSE",
    -- TX Initialization and Reset  
    TXPCSRESET_TIME                 => "00001",
    TXPMARESET_TIME                 => "00001",
    -- TX Receiver Detection        
    TX_RXDETECT_CFG                 => x"1832",
    TX_RXDETECT_REF                 => "100",
    -- JTAG                         
    ACJTAG_DEBUG_MODE               => '0',
    ACJTAG_MODE                     => '0',
    ACJTAG_RESET                    => '0',
    -- CDR                          
    CFOK_CFG                        => x"49000040E80",
    CFOK_CFG2                       => "0100000",
    CFOK_CFG3                       => "0100000",
    CFOK_CFG4                       => '0',
    CFOK_CFG5                       => x"0",
    CFOK_CFG6                       => "0000",
    RXOSCALRESET_TIME               => "00011",
    RXOSCALRESET_TIMEOUT            => "00000",
    -- PMA                          
    CLK_COMMON_SWING                => '0',
    RX_CLKMUX_EN                    => '1',
    TX_CLKMUX_EN                    => '1',
    ES_CLK_PHASE_SEL                => '0',
    USE_PCS_CLK_PHASE_SEL           => '0',
    PMA_RSV6                        => '0',
    PMA_RSV7                        => '0',
    -- TX Configuration Driver      
    TX_PREDRIVER_MODE               => '0',
    PMA_RSV5                        => '0',
    SATA_PLL_CFG                    => "VCO_3000MHZ",
    -- RX Fabric Clock Output Control
    RXOUT_DIV                       => 1, -- INFO: affects RXCDR_CFG attribute
    -- TX Fabric Clock Output Control
    TXOUT_DIV                       => 1, -- INFO: affects RXCDR_CFG attribute
    -- RX Phase Interpolator
    RXPI_CFG0                       => "000",
    RXPI_CFG1                       => '1',
    RXPI_CFG2                       => '1',
    -- RX Equalizer
    ADAPT_CFG0                      => x"00000",
    RXLPMRESET_TIME                 => "0001111",
    RXLPM_BIAS_STARTUP_DISABLE      => '0',
    RXLPM_CFG                       => "0110",
    RXLPM_CFG1                      => '0',
    RXLPM_CM_CFG                    => '0',
    RXLPM_GC_CFG                    => "111100010",
    RXLPM_GC_CFG2                   => "001",
    RXLPM_HF_CFG                    => "00001111110000",
    RXLPM_HF_CFG2                   => "01010",
    RXLPM_HF_CFG3                   => "0000",
    RXLPM_HOLD_DURING_EIDLE         => '0',
    RXLPM_INCM_CFG                  => '0',
    RXLPM_IPCM_CFG                  => '1',
    RXLPM_LF_CFG                    => "000000001111110000",
    RXLPM_LF_CFG2                   => "01010",
    RXLPM_OSINT_CFG                 => "100",
    -- TX Phase Interpolator PPM Controller
    TXPI_CFG0                       => "00",
    TXPI_CFG1                       => "00",
    TXPI_CFG2                       => "00",
    TXPI_CFG3                       => '0',
    TXPI_CFG4                       => '0',
    TXPI_CFG5                       => "000",
    TXPI_GREY_SEL                   => '0',
    TXPI_INVSTROBE_SEL              => '0',
    TXPI_PPMCLK_SEL                 => "TXUSRCLK2",
    TXPI_PPM_CFG                    => x"00",
    TXPI_SYNFREQ_PPM                => "001",
    -- Loopback
    LOOPBACK_CFG                    => '0',
    PMA_LOOPBACK_CFG                => '0',
    -- RX OOB Signalling
    RXOOB_CLK_CFG                   => "PMA",
    -- TX OOB Signalling
    TXOOB_CFG                       => '0',
    -- RX Buffer
    RXSYNC_MULTILANE                => '0',
    RXSYNC_OVRD                     => '0',
    RXSYNC_SKIP_DA                  => '0',
    -- TX Buffer
    TXSYNC_MULTILANE                => '0',
    TXSYNC_OVRD                     => '0',
    TXSYNC_SKIP_DA                  => '0'
  )
  port map
  (
    -- CPLL
    GTRSVD                          => "0000000000000000",
    PCSRSVDIN                       => "0000000000000000",
    TSTIN                           => "11111111111111111111",
    -- Dynamic Reconfiguration Port (DRP)
    DRPADDR                         => drp_addr,
    DRPCLK                          => ref_clk,
    DRPDI                           => drp_datain,
    DRPDO                           => drp_dataout,
    DRPEN                           => drp_en,
    DRPRDY                          => drp_rdy,
    DRPWE                           => drp_we,
    -- Clocking
    RXSYSCLKSEL                     => "00",   -- use PLL0 (hard coded)
    TXSYSCLKSEL                     => "00",   -- use PLL0 (hard coded)
    -- TX FPGA Interface Datapath Configuration
    TX8B10BEN                       => '1',
    -- GTPE2_CHANNEL Clocking
    PLL0CLK                         => pll0clk,
    PLL0REFCLK                      => pll0refclk,
    PLL1CLK                         => pll1clk,
    PLL1REFCLK                      => pll1refclk,
    -- Loopback
    LOOPBACK                        => loopen_i,
    -- PCI Express
    PHYSTATUS                       => open,
    RXRATE                          => "000",
    RXVALID                         => open,
    -- PMA Reserved
    PMARSVDIN3                      => '0',
    PMARSVDIN4                      => '0',
    -- Power-Down
    RXPD                            => "00",
    TXPD                            => "00",
    -- RX 8B/10B Decoder
    SETERRSTATUS                    => '0',
    -- RX Initialization and Reset
    EYESCANRESET                    => '0',
    RXUSERRDY                       => pll_lock,
    -- RX Margin Analysis
    EYESCANDATAERROR                => open,
    EYESCANMODE                     => '0',
    EYESCANTRIGGER                  => '0',
    -- RX Reset
    CLKRSVD0                        => '0',
    CLKRSVD1                        => '0',
    DMONFIFORESET                   => '0',
    DMONITORCLK                     => '0',
    RXPMARESETDONE                  => rx_pma_rst_done,
    SIGVALIDCLK                     => '0',
    -- RX CDR
    RXCDRFREQRESET                  => '0',
    RXCDRHOLD                       => '0',
    RXCDRLOCK                       => open,
    RXCDROVRDEN                     => '0',
    RXCDRRESET                      => '0',
    RXCDRRESETRSV                   => '0',
    RXOSCALRESET                    => '0',
    RXOSINTCFG                      => "0010",
    RXOSINTDONE                     => open,
    RXOSINTHOLD                     => '0',
    RXOSINTOVRDEN                   => '0',
    RXOSINTPD                       => '0',
    RXOSINTSTARTED                  => open,
    RXOSINTSTROBE                   => '0',
    RXOSINTSTROBESTARTED            => open,
    RXOSINTTESTOVRDEN               => '0',
    --RX Clock Correction
    RXCLKCORCNT                     => open,
    -- RX FPGA Interface Datapath Configuration
    RX8B10BEN                       => '1',
    -- RX FPGA Interface
    RXDATA                          => rx_data_full,
    RXUSRCLK                        => rx_clk,
    RXUSRCLK2                       => rx_clk,
    -- RX Pattern Checker
    RXPRBSERR                       => open,
    RXPRBSSEL                       => "000",
    RXPRBSCNTRESET                  => '0',
    -- RX 8B/10B Decoder
    RXCHARISCOMMA                   => open,
    RXCHARISK                       => rx_k_full,
    RXDISPERR                       => rx_disp_err,
    RXNOTINTABLE                    => rx_code_err,
    -- RX AFE
    GTPRXN                          => pad_rxn_i,
    GTPRXP                          => pad_rxp_i,
    PMARSVDIN2                      => '0',
    PMARSVDOUT0                     => open,
    PMARSVDOUT1                     => open,
    -- RX Buffer Bypass
    RXBUFRESET                      => '0',
    RXBUFSTATUS                     => rx_bufstatus,
    RXDDIEN                         => '0',
    RXDLYBYPASS                     => '1',
    RXDLYEN                         => '0',
    RXDLYOVRDEN                     => '0',
    RXDLYSRESET                     => '0',
    RXDLYSRESETDONE                 => open,
    RXPHALIGN                       => '0',
    RXPHALIGNDONE                   => open,
    RXPHALIGNEN                     => '0',
    RXPHDLYPD                       => '0',
    RXPHDLYRESET                    => '0',
    RXPHMONITOR                     => open,
    RXPHOVRDEN                      => '0',
    RXPHSLIPMONITOR                 => open,
    RXSTATUS                        => open,
    RXSYNCALLIN                     => '0',
    RXSYNCDONE                      => open,
    RXSYNCIN                        => '0',
    RXSYNCMODE                      => '0',
    RXSYNCOUT                       => open,
    -- RX Byte and Word Alignment
    RXBYTEISALIGNED                 => rx_synced_o,
    RXBYTEREALIGN                   => open,
    RXCOMMADET                      => open,
    RXCOMMADETEN                    => '1',
    RXMCOMMAALIGNEN                 => rx_resync_i,
    RXPCOMMAALIGNEN                 => rx_resync_i,
    RXSLIDE                         => '0',
    -- RX Channel Bonding
    RXCHANBONDSEQ                   => open,
    RXCHBONDEN                      => '0',
    RXCHBONDI                       => "0000",
    RXCHBONDLEVEL                   => "000",
    RXCHBONDMASTER                  => '0',
    RXCHBONDO                       => open,
    RXCHBONDSLAVE                   => '0',
    -- RX Channel Bonding
    RXCHANISALIGNED                 => open,
    RXCHANREALIGN                   => open,
    -- RX Decision Feedback Equalizer (DFE)
    DMONITOROUT                     => open,
    RXADAPTSELTEST                  => "00000000000000",
    RXDFEXYDEN                      => '0',
    RXOSINTEN                       => '1',
    RXOSINTID0                      => "0000",
    RXOSINTNTRLEN                   => '0',
    RXOSINTSTROBEDONE               => open,
    -- RX Driver, OOB Signalling, Coupling and Equalizer, CDR
    RXLPMLFOVRDEN                   => '0',
    RXLPMOSINTNTRLEN                => '0',
    -- RX Equalizer
    RXLPMHFHOLD                     => '0',
    RXLPMHFOVRDEN                   => '0',
    RXLPMLFHOLD                     => '0',
    RXOSHOLD                        => '0',
    RXOSOVRDEN                      => '0',
    -- RX Fabric ClocK Output Control
    RXRATEDONE                      => open,
    RXRATEMODE                      => '0',
    RXOUTCLK                        => open,
    RXOUTCLKFABRIC                  => open,
    RXOUTCLKPCS                     => open,
    RXOUTCLKSEL                     => "010",
    -- RX Gearbox
    RXDATAVALID                     => open,
    RXHEADER                        => open,
    RXHEADERVALID                   => open,
    RXSTARTOFSEQ                    => open,
    RXGEARBOXSLIP                   => '0',
    -- RX Initialization and Reset
    GTRXRESET                       => rx_rst_seqout,
    RXLPMRESET                      => '0',
    RXOOBRESET                      => '0',
    RXPCSRESET                      => '0',
    RXPMARESET                      => '0',
    -- RX OOB Signalling
    RXCOMSASDET                     => open,
    RXCOMWAKEDET                    => open,
    RXCOMINITDET                    => open,
    RXELECIDLE                      => open,
    RXELECIDLEMODE                  => "11",
    -- RX Polarity Control
    RXPOLARITY                      => '0',
    -- RX Initialization and Reset
    RXRESETDONE                     => rx_rst_done,
    -- TX Buffer Bypass
    TXPHDLYTSTCLK                   => '0',
    -- TX Configurable Driver
    TXPOSTCURSOR                    => "00000",
    TXPOSTCURSORINV                 => '0',
    TXPRECURSOR                     => "00000",
    TXPRECURSORINV                  => '0',
    -- TX Fabric Clock Output Control
    TXRATEMODE                      => '0',
    -- TX Initialization and Reset
    CFGRESET                        => '0',
    GTTXRESET                       => tx_rst,
    PCSRSVDOUT                      => open,
    TXUSERRDY                       => pll_lock,
    -- TX Phase Interpolator PPM Controller
    TXPIPPMEN                       => '0',
    TXPIPPMOVRDEN                   => '0',
    TXPIPPMPD                       => '0',
    TXPIPPMSEL                      => '1',
    TXPIPPMSTEPSIZE                 => "00000",
    -- Transceiver Reset Mode Operation
    GTRESETSEL                      => '0',
    RESETOVRD                       => '0',
    -- TX Reset
    TXPMARESETDONE                  => tx_pma_rst_done,
    -- TX Configurable Driver
    PMARSVDIN0                      => '0',
    PMARSVDIN1                      => '0',
    -- TX FPGA Interface
    TXDATA                          => tx_data_full,
    TXUSRCLK                        => tx_clk,
    TXUSRCLK2                       => tx_clk,
    -- TX PCI Express
    TXELECIDLE                      => '0',
    TXMARGIN                        => "000",
    TXRATE                          => "000",
    TXSWING                         => '0',
    -- TX Pattern Generator
    TXPRBSFORCEERR                  => '0',
    -- TX 8B/10B Encoder
    TX8B10BBYPASS                   => "0000",
    TXCHARDISPMODE                  => "0000",
    TXCHARDISPVAL                   => "0000",
    TXCHARISK(3 downto 2)           => "00",
    TXCHARISK(1 downto 0)           => tx_k_i,
    -- TX Buffer Bypass
    TXDLYBYPASS                     => '1',
    TXDLYEN                         => '0',
    TXDLYHOLD                       => '0',
    TXDLYOVRDEN                     => '0',
    TXDLYSRESET                     => '0',
    TXDLYSRESETDONE                 => open,
    TXDLYUPDOWN                     => '0',
    TXPHALIGN                       => '0',
    TXPHALIGNDONE                   => open,
    TXPHALIGNEN                     => '0',
    TXPHDLYPD                       => '0',
    TXPHDLYRESET                    => '0',
    TXPHINIT                        => '0',
    TXPHINITDONE                    => open,
    TXPHOVRDEN                      => '0',
    -- TX Buffer
    TXBUFSTATUS                     => open,
    -- TX Buffer and Phase Alignment
    TXSYNCALLIN                     => '0',
    TXSYNCDONE                      => open,
    TXSYNCIN                        => '0',
    TXSYNCMODE                      => '0',
    TXSYNCOUT                       => open,
    -- TX Configurable Driver
    GTPTXN                          => pad_txn_o,
    GTPTXP                          => pad_txp_o,
    TXBUFDIFFCTRL                   => "100",
    TXDEEMPH                        => '0',
    TXDIFFCTRL                      => "1000",
    TXDIFFPD                        => '0',
    TXINHIBIT                       => '0',
    TXMAINCURSOR                    => "0000000",
    TXPISOPD                        => '0',
    -- TX Fabric Clock Output Control
    TXOUTCLK                        => tx_clk_bufin,
    TXOUTCLKFABRIC                  => open,
    TXOUTCLKPCS                     => open,
    TXOUTCLKSEL                     => "010",
    TXRATEDONE                      => open,
    -- TX Gearbox
    TXGEARBOXREADY                  => open,
    TXHEADER                        => "000",
    TXSEQUENCE                      => "0000000",
    TXSTARTSEQ                      => '0',
    -- TX Initialization and Reset
    TXPCSRESET                      => '0',
    TXPMARESET                      => '0',
    TXRESETDONE                     => tx_rst_done,
    -- TX OOB Signalling
    TXCOMFINISH                     => open,
    TXCOMINIT                       => '0',
    TXCOMSAS                        => '0',
    TXCOMWAKE                       => '0',
    TXPDELECIDLEMODE                => '0',
    -- TX Polarity Control
    TXPOLARITY                      => '0',
    -- TX Receiver Detection
    TXDETECTRX                      => '0',
    -- TX Pattern Generator
    TXPRBSSEL                       => "000"
  );

  -- GTP reset sequence upon FPGA configuration (AR# 53561)
  -- Based on code generated by Vivado GT wizard (<gtname>_gtrxreset_seq.vhd)
  -- TODO: replace sync_block by gc_sync_ffs
  gen_gtrxreset_seq : if g_SIMULATION /= "TRUE" generate
    cmp_gtrxreset_seq_0 : gtrxreset_seq
    port map
    (
      RST             =>  rst_synced,
      GTRXRESET_IN    =>  rx_rst,
      RXPMARESETDONE  =>  rx_pma_rst_done,
      GTRXRESET_OUT   =>  rx_rst_seqout,
      DRP_OP_DONE     =>  drp_done,
      DRPCLK          =>  ref_clk,
      DRPEN           =>  drp_en,
      DRPADDR         =>  drp_addr,
      DRPWE           =>  drp_we,
      DRPDO           =>  drp_dataout,
      DRPDI           =>  drp_datain,
      DRPRDY          =>  drp_rdy
    );
  end generate;

  gen_gtrxreset_seq_sim : if g_SIMULATION = "TRUE" generate
    cmp_gtrxreset_seq_0 : gtrxreset_seq_sim
    port map
    (
      RST             =>  rst_synced,
      GTRXRESET_IN    =>  rx_rst,
      RXPMARESETDONE  =>  rx_pma_rst_done,
      GTRXRESET_OUT   =>  rx_rst_seqout,
      DRP_OP_DONE     =>  drp_done,
      DRPCLK          =>  ref_clk,
      DRPEN           =>  drp_en,
      DRPADDR         =>  drp_addr,
      DRPWE           =>  drp_we,
      DRPDO           =>  drp_dataout,
      DRPDI           =>  drp_datain,
      DRPRDY          =>  drp_rdy
    );
  end generate;

  -- Quad GTP PLL instance
  cmp_gtpll : GTPE2_COMMON
  generic map
  (
    -- Simulation
    SIM_RESET_SPEEDUP       => g_SIMULATION,
    SIM_PLL0REFCLK_SEL      => "001",
    SIM_PLL1REFCLK_SEL      => "001",
    SIM_VERSION             => "2.0",
    -- PLL Dividers
    PLL0_FBDIV              => c_PLLFBDIV,
    PLL0_FBDIV_45           => c_PLLFBDIV45,
    PLL0_REFCLK_DIV         => c_PLLREFDIV,
    PLL1_FBDIV              => 1,
    PLL1_FBDIV_45           => 4,
    PLL1_REFCLK_DIV         => 1,
    -- Common Block
    BIAS_CFG                => x"0000000000050001",
    COMMON_CFG              => x"00000000",
    -- PLL
    PLL0_CFG                => x"01F03DC",
    PLL0_DMON_CFG           => '0',
    PLL0_INIT_CFG           => x"00001E",
    PLL0_LOCK_CFG           => x"1E8",
    PLL1_CFG                => x"01F03DC",
    PLL1_DMON_CFG           => '0',
    PLL1_INIT_CFG           => x"00001E",
    PLL1_LOCK_CFG           => x"1E8",
    PLL_CLKOUT_CFG          => x"00",
    -- Reserved
    RSVD_ATTR0              => x"0000",
    RSVD_ATTR1              => x"0000"
  )
  port map
  (
    DMONITOROUT             => open,
    -- Dynamic Reconfiguration Port (DRP)
    DRPADDR                 => "00000000",
    DRPCLK                  => '0',
    DRPDI                   => "0000000000000000",
    DRPDO                   => open,
    DRPEN                   => '0',
    DRPRDY                  => open,
    DRPWE                   => '0',
    -- GTPE2_COMMON Clocking
    GTGREFCLK0              => '0',
    GTGREFCLK1              => '0',
    GTEASTREFCLK0           => gteastrefclk0,
    GTEASTREFCLK1           => gteastrefclk1,
    GTREFCLK0               => gtrefclk0,
    GTREFCLK1               => gtrefclk1,
    GTWESTREFCLK0           => gtwestrefclk0,
    GTWESTREFCLK1           => gtwestrefclk1,
    PLL0OUTCLK              => pll0clk,
    PLL0OUTREFCLK           => pll0refclk,
    PLL1OUTCLK              => pll1clk,
    PLL1OUTREFCLK           => pll1refclk,
    -- PLL                  
    PLL0FBCLKLOST           => open,
    PLL0LOCK                => pll_lock,
    PLL0LOCKDETCLK          => '0',
    PLL0LOCKEN              => '1',
    PLL0PD                  => '0',
    PLL0REFCLKLOST          => open,
    PLL0REFCLKSEL           => pll0refclksel,
    PLL0RESET               => pll_rst,
    PLL1FBCLKLOST           => open,
    PLL1LOCK                => open,
    PLL1LOCKDETCLK          => '0',
    PLL1LOCKEN              => '1',
    PLL1PD                  => '1',
    PLL1REFCLKLOST          => open,
    PLL1REFCLKSEL           => "001",
    PLL1RESET               => '0',
    -- Common Block         
    BGRCALOVRDENB           => '1',
    PLLRSVD1                => "0000000000000000",
    PLLRSVD2                => "00000",
    REFCLKOUTMONITOR0       => open,
    REFCLKOUTMONITOR1       => open,
    -- RX AFE               
    PMARSVDOUT              => open,
    -- QPLL                 
    BGBYPASSB               => '1',
    BGMONITORENB            => '1',
    BGPDB                   => '1',
    BGRCALOVRD              => "11111",
    PMARSVD                 => "00000000",
    RCALENB                 => '1'
  );

  -- GT reference clock input buffer
  gen_refclk_ibufbds : if g_REFCLK = "REFCLK0" or g_REFCLK = "REFCLK1" generate
    cmp_ibufbds_gte2 : IBUFDS_GTE2
    port map
    (
      O       => ref_clk,
      ODIV2   => open,
      CEB     => '0',
      I       => pad_refclkp_i,
      IB      => pad_refclkn_i
    );
  end generate;

  gen_refclk0 : if g_REFCLK = "REFCLK0" generate
    gtrefclk0     <= ref_clk;
    gtrefclk1     <= '0';
    gteastrefclk0 <= '0';
    gteastrefclk1 <= '0';
    gtwestrefclk0 <= '0';
    gtwestrefclk1 <= '0';
    pll0refclksel <= "001";
  end generate;

  gen_refclk1 : if g_REFCLK = "REFCLK1" generate
    gtrefclk0     <= '0';
    gtrefclk1     <= ref_clk;
    gteastrefclk0 <= '0';
    gteastrefclk1 <= '0';
    gtwestrefclk0 <= '0';
    gtwestrefclk1 <= '0';
    pll0refclksel <= "010";    
  end generate;

  gen_eastrefclk0 : if g_REFCLK = "EASTREFCLK0" generate
    gtrefclk0     <= '0';
    gtrefclk1     <= '0';
    gteastrefclk0 <= ref_clk;
    gteastrefclk1 <= '0';
    gtwestrefclk0 <= '0';
    gtwestrefclk1 <= '0';
    pll0refclksel <= "011";
  end generate;

  gen_eastrefclk1 : if g_REFCLK = "EASTREFCLK1" generate
    gtrefclk0     <= '0';
    gtrefclk1     <= '0';
    gteastrefclk0 <= '0';
    gteastrefclk1 <= ref_clk;
    gtwestrefclk0 <= '0';
    gtwestrefclk1 <= '0';
    pll0refclksel <= "100";
  end generate;

  gen_gtwestrefclk0 : if g_REFCLK = "WESTREFCLK0" generate
    gtrefclk0     <= '0';
    gtrefclk1     <= '0';
    gteastrefclk0 <= '0';
    gteastrefclk1 <= '0';
    gtwestrefclk0 <= ref_clk;
    gtwestrefclk1 <= '0';
    pll0refclksel <= "101";
  end generate;

  gen_gtwestrefclk1 : if g_REFCLK = "WESTREFCLK1" generate
    gtrefclk0     <= '0';
    gtrefclk1     <= '0';
    gteastrefclk0 <= '0';
    gteastrefclk1 <= '0';
    gtwestrefclk0 <= '0';
    gtwestrefclk1 <= ref_clk;
    pll0refclksel <= "110";
  end generate;

  -- User clock global buffer
  cmp_tx_clk_bufg : BUFG
  port map
  (
    I => tx_clk_bufin,
    O => tx_clk
  );

  tx_clk_o      <= tx_clk;

  -- When RX elastic buffer is in use RXUSRCLK is driven by TXOUTCLK
  rx_clk        <= tx_clk;
  rx_clk_o      <= rx_clk;

  -- RX outputs
  rx_data_o     <= rx_data_full(15 downto 0);
  rx_k_o        <= rx_k_full(1 downto 0);
  rx_enc_err_o  <= rx_disp_err(1) or rx_disp_err(0) or rx_code_err(1) or rx_code_err(0);
  rx_buf_err_o  <= rx_bufstatus(2);

  -- TX input: pad unused data bits
  tx_data_full  <= "0000000000000000" & tx_data_i;

  -- RX reset and ready
  rx_rst        <= not pll_rst and (not pll_lock or rx_rst_i);
  rx_rdy_o      <= pll_lock and tx_rst_done and rx_rst_done;

  -- TX reset and ready
  tx_rst        <= not pll_rst and (not pll_lock or tx_rst_i);
  tx_rdy_o      <= pll_lock and tx_rst_done;

  -- Detect edge and synchronize with GT reference clock
  cmp_rst_sync : gc_sync_ffs
  generic map
  (
    g_sync_edge => "positive"
  )
  port map
  (
    clk_i       => ref_clk,
    rst_n_i     => '1',
    data_i      => rst_i,
    ppulse_o    => rst_synced
  );

  -- Wait a minimum of 500 ns after configuration is complete as per UG482
  -- "GTP Transceiver TX/RX Reset in Response to Completion of Configuration"
  p_rst_wait : process(ref_clk, rst_synced) is
    variable reset_cnt : integer range 0 to c_RST_DELAY := 0;
  begin
    if rst_synced = '1' then
      reset_cnt := 0;
      pll_rst <= '1';
    elsif rising_edge(ref_clk) then
      if reset_cnt = c_RST_DELAY then
        pll_rst <= '0';
      else
        reset_cnt := reset_cnt + 1;
        pll_rst <= '1';
      end if;
    end if;
  end process;

end rtl;
